// $Id: $
// File name:   tb_sha256_640.sv
// Created:     11/1/2014
// Author:      Kyle Chynoweth
// Lab Section: 01
// Version:     1.0  Initial Design Entry
// Description: SHA256 80-octet test bench
module tb_sha256_640();
endmodule