// $Id: $
// File name:   hmac_sha256_32.sv
// Created:     11/15/2014
// Author:      Kyle Chynoweth
// Lab Section: 01
// Version:     1.0  Initial Design Entry
// Description: Common module for all hmac_sha256_x blocks
